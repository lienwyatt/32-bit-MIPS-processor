---------------------------------------------------------------------------------
-- Memory unit
-- contains all memory for the a 32 bit MIPS processor
-- includes data memory which can be read and written to as well as read only 
-- instruction memory
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity memory_unit is
port
(
ab1: in std_logic_vector(31 downto 0); -- pc (address of instruction)
ib1: out std_logic_vector(31 downto 0); -- instruction fetched from memory

ab2: in std_logic_vector(31 downto 0); --  address of data (to be fetched or written to)
db2: in std_logic_vector(31 downto 0); -- carries the data to be written to memory
write_en : in std_logic; -- write enable
db3: out std_logic_vector(31 downto 0); -- data out

clear: in std_logic; -- clear bit (for data memory)
clock : in std_logic; -- clock signal
switches:in std_logic_vector(15 downto 0)
);
end memory_unit;

architecture Behavioral of memory_unit is

signal inst_addr : std_logic_vector(31 downto 0);
signal inst : std_logic_vector(31 downto 0); -- instruction that'll go out on ib1

signal data_addr : std_logic_vector(31 downto 0);
signal data_in : std_logic_vector(31 downto 0);
signal data_out : std_logic_vector(31 downto 0);


-- size of memory is 64x32 (64 32-bit locations)
type rom is array (0 to 63) of std_logic_vector(31 downto 0);
type ram is array (0 to 63) of std_logic_vector(31 downto 0);

--instruction memory
--instruction memory (count instances progeam). Remove spaces before implementing. They are for documentation/debug purposes
constant inst_mem : rom :=
(  
"10001100000000100000000000011100","00000000000000000011000000100000","00000000000000000001100000100000","00100100000001000000000000010101",--lw, add, add, addi, 
"10001100011001010000000000000000", --load
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000",  
"00100000011000110000000000000001","00010000101000100000000000001111", --branch
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"00010100011001000000000000001011",--instruction 60(decimal) branch
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000",  
"00001000000000000000000000011111", --instruction 80(decimal) jump
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000",
"00000000110000010011000000100000","00001000000000000000000000000100",--instruction 104 jump
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000",
"10101100000001100000000000011111",  
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"00001000000000000000000000101000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", --jump for infintite loop of noops
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000",
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000", 
"11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000","11111100000000000000000000000000"
--"11111100000000000000000000000000", "11111100000000000000000000000000", "11111100000000000000000000000000", "11111100000000000000000000000000",
--"11111100000000000000000000000000" "11111100000000000000000000000000", "11111100000000000000000000000000", "11111100000000000000000000000000"
--"11111100000000000000000000000000", "11111100000000000000000000000000", "11111100000000000000000000000000", "11111100000000000000000000000000", 
);

--DATA Memory. In this example the array is searched for "110" or 6, the destination is on line 31, location 0x20. It should find 3 instances.
signal data_mem : ram := 
(
--"00000000000000000000000000000001", "00000000000000000000000000001100", "00000000000000000000000000000110", "00000000000000000000000000000110", 
--"00000000000000000000000000000001", "00000000000000000000000000000110", "00000000000000000000000000000001", "00000000000000000000000000000101", 
--"00000000000000000000000000001111", "00000000000000000000000000000011", "00000000000000000000000000000001", "00000000000000000000000000000011", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000111", "00000000000000000000000000000001", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000100", "00000000000000000000000000000000", "00000000000000000000000000000001", 
--"00000000000000000000000000000110", "00000000000000000000000000001000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000"


"00000000000000000000000000000001", "00000000000000000000000000001100", "00000000000000000000000000000110", "00000000000000000000000000000110", 
"00000000000000000000000000000001", "00000000000000000000000000000110", "00000000000000000000000000000001", "00000000000000000000000000000101", 
"00000000000000000000000000001111", "00000000000000000000000000000011", "00000000000000000000000000000001", "00000000000000000000000000000011", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"00000000000000000000000000000111", "00000000000000000000000000000001", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"00000000000000000000000000000110", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", 
"10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000", "10000000000000000000000000000000"

);

--data memory
signal data_mem_cleared : ram := 
(

"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", 
"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000" 
);


begin

inst_addr <= ab1;
data_addr <= ab2;
data_in <= db2;

-- process to get next instruction
process(clock)
begin
	if(clock = '1' and clock' event) then
		inst <= inst_mem(to_integer(unsigned(inst_addr))/4);
	end if;
end process;
data_out <= data_mem(to_integer(unsigned(data_addr))); -- read data CHANGE THISSSSS


--process to read/write data, data memory can be cleared as well
process(clock, clear)
begin
	if(clear = '1') then
		if (clock' event and clock='1') then
			data_mem(28)<="0000000000000000" & switches;
		END IF;
	else
		if(clock = '1' and clock' event) then
			-- write data to memory
			if(write_en = '1') then
				data_mem(to_integer(unsigned(data_addr))) <= data_in;
			end if;
		end if;
	end if;
end process;

ib1 <= inst;
db3 <= data_out;


end Behavioral;
